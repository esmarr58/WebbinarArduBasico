module S1L1
	 (
		input 	A,
		input 	B,
		output   Y
	 );
        assign Y = A & B;
    endmodule